,topic_name,topic_details,topic_url
0,3D,3D modeling is the process of virtually developing the surface and structure of a 3D object.,https://github.com/topics/3d
1,Ajax,Ajax is a technique for creating interactive web applications.,https://github.com/topics/ajax
2,Algorithm,Algorithms are self-contained sequences that carry out a variety of tasks.,https://github.com/topics/algorithm
3,Amp,Amp is a non-blocking concurrency library for PHP.,https://github.com/topics/amphp
4,Android,Android is an operating system built by Google designed for mobile devices.,https://github.com/topics/android
5,Angular,Angular is an open source web application platform.,https://github.com/topics/angular
6,Ansible,Ansible is a simple and powerful automation engine.,https://github.com/topics/ansible
7,API,An API (Application Programming Interface) is a collection of protocols and subroutines for building software.,https://github.com/topics/api
8,Arduino,Arduino is an open source hardware and software company and maker community.,https://github.com/topics/arduino
9,ASP.NET,ASP.NET is a web framework for building modern web apps and services.,https://github.com/topics/aspnet
10,Atom,Atom is a open source text editor built with web technologies.,https://github.com/topics/atom
11,Awesome Lists,An awesome list is a list of awesome things curated by the community.,https://github.com/topics/awesome
12,Amazon Web Services,Amazon Web Services provides on-demand cloud computing platforms on a subscription basis.,https://github.com/topics/aws
13,Azure,Azure is a cloud computing service created by Microsoft.,https://github.com/topics/azure
14,Babel,"Babel is a compiler for writing next generation JavaScript, today.",https://github.com/topics/babel
15,Bash,Bash is a shell and command language interpreter for the GNU operating system.,https://github.com/topics/bash
16,Bitcoin,Bitcoin is a cryptocurrency developed by Satoshi Nakamoto.,https://github.com/topics/bitcoin
17,Bootstrap,"Bootstrap is an HTML, CSS, and JavaScript framework.",https://github.com/topics/bootstrap
18,Bot,A bot is an application that runs automated tasks over the Internet.,https://github.com/topics/bot
19,C,C is a general purpose programming language that first appeared in 1972.,https://github.com/topics/c
20,Chrome,Chrome is a web browser from the tech company Google.,https://github.com/topics/chrome
21,Chrome extension,Google Chrome Extensions are add-ons that allow users to customize their Chrome web browser.,https://github.com/topics/chrome-extension
22,Command line interface,"A CLI, or command-line interface, is a console that helps users issue commands to a program.",https://github.com/topics/cli
23,Clojure,"Clojure is a dynamic, general-purpose programming language.",https://github.com/topics/clojure
24,Code quality,"Automate your code review with style, quality, security, and testâ€‘coverage checks when you need them.",https://github.com/topics/code-quality
25,Code review,Ensure your code meets quality standards and ship with confidence.,https://github.com/topics/code-review
26,Compiler,Compilers are software that translate higher-level programming languages to lower-level languages (e.g. machine code).,https://github.com/topics/compiler
27,Continuous integration,"Automatically build and test your code as you push it upstream, preventing bugs from being deployed to production.",https://github.com/topics/continuous-integration
28,COVID-19,The coronavirus disease 2019 (COVID-19) is an infectious disease caused by SARS-CoV-2.,https://github.com/topics/covid-19
29,C++,C++ is a general purpose and object-oriented programming language.,https://github.com/topics/cpp
